/******************************************************************************

SDRAM ctrl

******************************************************************************/

module sdram_ctrl
(
    input clk,
    input clk_shift,
    input rst_n
);

endmodule
